library verilog;
use verilog.vl_types.all;
entity memory_test_vlg_vec_tst is
end memory_test_vlg_vec_tst;
