library verilog;
use verilog.vl_types.all;
entity decoBCD_vlg_vec_tst is
end decoBCD_vlg_vec_tst;
